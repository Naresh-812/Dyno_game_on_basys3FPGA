module line_rom(vc,outl);
input [10:0]vc;
output reg[699:0]outl;
always@(vc)
begin
case(vc-10'd400)
4'd0:outl<=700'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
4'd1:outl<=700'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
4'd2:outl<=700'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
4'd3:outl<=700'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
4'd4:outl<=700'b000011111000000000001111100000000000000001111100000000000000000000011111000000000000001111100000000000111110000000000000001111100000000000000000011111000000000000000000011111000000000001111100000000000011111000000000000000011111000000000000000000000111110000000000000000011111000000000000000111110000000000000000111110000000000000000001111100000000000001111100000000000000011111000000000000000000001111100000000000000000000000111110000000000000000000000111110000000000000011111000000000000000000001111100000000000000011111000000000000000000000011111000000000000000000001111100000000000000111110000000000000000000011111000000000000000000111110000000000000011111000000000000011111000000000001111100000;
4'd5:outl<=700'b000011111000000000001111100000000000000001111100000000000000000000011111000000000000001111100000000000111110000000000000001111100000000000000000011111000000000000000000011111000000000001111100000000000011111000000000000000011111000000000000000000000111110000000000000000011111000000000000000111110000000000000000111110000000000000000001111100000000000001111100000000000000011111000000000000000000001111100000000000000000000000111110000000000000000000000111110000000000000011111000000000000000000001111100000000000000011111000000000000000000000011111000000000000000000001111100000000000000111110000000000000000000011111000000000000000000111110000000000000011111000000000000011111000000000001111100000;
4'd6:outl<=700'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
4'd7:outl<=700'b000000000000001111100000000000111110000000000000000111110000000000000000000001111100000000000000111110000000000011111000000000000000111110000000000000000001111100000000000000000001111100000000000111110000000000001111100000000000000001111100000000000000000000011111000000000000000001111100000000000000011111000000000000000011111000000000000000000111110000000000000111110000000000000001111100000000000000000000111110000000000000000000000011111000000000000000000000011111000000000000001111100000000000000000000111110000000000000001111100000000000000000000001111100000000000000000000111110000000000000011111000000000000000000001111100000000000000000011111000000000000001111100000000000001111100000000000;
4'd8:outl<=700'b000000000000001111100000000000111110000000000000000111110000000000000000000001111100000000000000111110000000000011111000000000000000111110000000000000000001111100000000000000000001111100000000000111110000000000001111100000000000000001111100000000000000000000011111000000000000000001111100000000000000011111000000000000000011111000000000000000000111110000000000000111110000000000000001111100000000000000000000111110000000000000000000000011111000000000000000000000011111000000000000001111100000000000000000000111110000000000000001111100000000000000000000001111100000000000000000000111110000000000000011111000000000000000000001111100000000000000000011111000000000000001111100000000000001111100000000000;
4'd9:outl<=700'b000000000000001111100000000000111110000000000000000111110000000000000000000001111100000000000000111110000000000011111000000000000000111110000000000000000001111100000000000000000001111100000000000111110000000000001111100000000000000001111100000000000000000000011111000000000000000001111100000000000000011111000000000000000011111000000000000000000111110000000000000111110000000000000001111100000000000000000000111110000000000000000000000011111000000000000000000000011111000000000000001111100000000000000000000111110000000000000001111100000000000000000000001111100000000000000000000111110000000000000011111000000000000000000001111100000000000000000011111000000000000001111100000000000001111100000000000;
endcase
end
endmodule