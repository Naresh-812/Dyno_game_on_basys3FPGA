module dino_rom(clk,addr_dino,outd);
input clk;
input [11:0]addr_dino;
output reg [21:0] outd;

always @(posedge clk)
begin
case(addr_dino)
//////////////////////////////////////////////////////////////////////////
12'h000:outd<=22'b0000000000000000000000;
12'h001:outd<=22'b0000000000000000000000;
12'h002:outd<=22'b0011111111000000000000;
12'h003:outd<=22'b0011111111000000000000;
12'h004:outd<=22'b0111111111100000000000;
12'h005:outd<=22'b0111111101100000000000;
12'h006:outd<=22'b0111111101100000000000;
12'h007:outd<=22'b0111111111100000000000;
12'h008:outd<=22'b0111111111100000000000;
12'h009:outd<=22'b0111111111100000000000;
12'h00a:outd<=22'b0111111111100000000000;
12'h00b:outd<=22'b0111111111100000000000;
12'h00c:outd<=22'b0111111111100000000000;
12'h00d:outd<=22'b0000001111100000000000;
12'h00e:outd<=22'b0000001111100000000000;
12'h00f:outd<=22'b0001111111100000000000;
12'h010:outd<=22'b0001111111100000000000;
12'h011:outd<=22'b0000000111110000000010;
12'h012:outd<=22'b0000000111110000000010;
12'h013:outd<=22'b0000000111111000000010;
12'h014:outd<=22'b0000000111111000000010;
12'h015:outd<=22'b0000011111111110000110;
12'h016:outd<=22'b0000011111111110000110;
12'h017:outd<=22'b0000010111111111001110;
12'h018:outd<=22'b0000010111111111001110;
12'h019:outd<=22'b0000000111111111111110;
12'h01a:outd<=22'b0000000111111111111110;
12'h01b:outd<=22'b0000000111111111111110;
12'h01c:outd<=22'b0000000111111111111110;
12'h01d:outd<=22'b0000000111111111111100;
12'h01e:outd<=22'b0000000011111111111100;
12'h01f:outd<=22'b0000000011111111111000;
12'h020:outd<=22'b0000000011111111111000;
12'h021:outd<=22'b0000000001111111110000;
12'h022:outd<=22'b0000000001111111110000;
12'h023:outd<=22'b0000000000111111100000;
12'h024:outd<=22'b0000000000111111100000;
12'h025:outd<=22'b0000000000110011000000;
12'h026:outd<=22'b0000000000110011000000;
12'h027:outd<=22'b0000000000100110000000;
12'h028:outd<=22'b0000000000100110000000;
12'h029:outd<=22'b0000000000100000000000;
12'h02a:outd<=22'b0000000000100000000000;
12'h02b:outd<=22'b0000000001100000000000;
12'h02c:outd<=22'b0000000001100000000000;
12'h02d:outd<=22'b0000000000000000000000;
12'h02e:outd<=22'b0000000000000000000000;

///////////////////////////////////////////////////////////////////////////////////////////

12'h100:outd<=22'b0000000000000000000000;
12'h101:outd<=22'b0000000000000000000000;
12'h102:outd<=22'b0011111111000000000000;
12'h103:outd<=22'b0011111111000000000000;
12'h104:outd<=22'b0111111111100000000000;
12'h105:outd<=22'b0111111101100000000000;
12'h106:outd<=22'b0111111101100000000000;
12'h107:outd<=22'b0111111111100000000000;
12'h108:outd<=22'b0111111111100000000000;
12'h109:outd<=22'b0111111111100000000000; 
12'h10a:outd<=22'b0111111111100000000000;
12'h10b:outd<=22'b0111111111100000000000;
12'h10c:outd<=22'b0111111111100000000000;
12'h10d:outd<=22'b0000001111100000000000;
12'h10e:outd<=22'b0000001111100000000000;
12'h10f:outd<=22'b0001111111100000000000;
12'h110:outd<=22'b0001111111100000000000;
12'h111:outd<=22'b0000000111110000000010;
12'h112:outd<=22'b0000000111110000000010;
12'h113:outd<=22'b0000000111111000000010;
12'h114:outd<=22'b0000000111111000000010;
12'h115:outd<=22'b0000011111111110000110;
12'h116:outd<=22'b0000011111111110000110;
12'h117:outd<=22'b0000010111111111001110;
12'h118:outd<=22'b0000010111111111001110;
12'h119:outd<=22'b0000000111111111111110;
12'h11a:outd<=22'b0000000111111111111110;
12'h11b:outd<=22'b0000000111111111111110;
12'h11c:outd<=22'b0000000111111111111110;
12'h11d:outd<=22'b0000000111111111111100;
12'h11e:outd<=22'b0000000011111111111100;
12'h12f:outd<=22'b0000000011111111111000;
12'h120:outd<=22'b0000000011111111111000;
12'h121:outd<=22'b0000000001111111110000;
12'h122:outd<=22'b0000000001111111110000;
12'h123:outd<=22'b0000000000111111100000;
12'h124:outd<=22'b0000000000111111100000;
12'h125:outd<=22'b0000000001100111000000;
12'h126:outd<=22'b0000000001100111000000;
12'h127:outd<=22'b0000000000000011000000;
12'h128:outd<=22'b0000000000000011000000;
12'h129:outd<=22'b0000000000000001000000;
12'h12a:outd<=22'b0000000000000001000000;
12'h12b:outd<=22'b0000000000000011000000;
12'h12c:outd<=22'b0000000000000011000000;
12'h12d:outd<=22'b0000000000000000000000;
12'h12e:outd<=22'b0000000000000000000000;   
        endcase
    end
endmodule

