module bird_rom(addrb,outb);
input [11:0]addrb;
output reg [49:0]outb;
always@(addrb)
begin
case(addrb)
12'h000:outb<=50'b00000000000000000000000000000000000000000000000000;
12'h001:outb<=50'b00000000000000000000001100000000000000000000000000;
12'h002:outb<=50'b00000000000000000000001100000000000000000000000000;
12'h003:outb<=50'b00000000000000000000001111000000000000000000000000;
12'h004:outb<=50'b00000000000000000000001111000000000000000000000000;
12'h005:outb<=50'b00000000000000000000001111110000000000000000000000;
12'h006:outb<=50'b00000000000000000000001111110000000000000000000000;
12'h007:outb<=50'b00000000000000000000001111111100000000000000000000;
12'h008:outb<=50'b00000000000000000000001111111100000000000000000000;
12'h009:outb<=50'b00000000000000000000001111111100000000000000000000;
12'h00a:outb<=50'b00000000000000000000001111111100000000000000000000;
12'h00b:outb<=50'b00000000000011110000001111111111000000000000000000;
12'h00c:outb<=50'b00000000000011110000001111111111000000000000000000;
12'h00d:outb<=50'b00000000001111111100001111111111110000000000000000;
12'h00e:outb<=50'b00000000001111111100001111111111110000000000000000;
12'h00f:outb<=50'b00000000111111111111001111111111111100000000000000;
12'h010:outb<=50'b00000001111111111111001111111111111100000000000000;
12'h011:outb<=50'b00000011111111111111001111111111111111000000000000;
12'h012:outb<=50'b00000111111111111111001111111111111111000000000000;
12'h013:outb<=50'b00001111111111111111111111111111111111111111110000;
12'h014:outb<=50'b00001111111111111111111111111111111111111111110000;
12'h015:outb<=50'b00000000000000001111111111111111111111110000000000;
12'h016:outb<=50'b00000000000000001111111111111111111111110000000000;
12'h017:outb<=50'b00000000000000000000111111111111111111111111000000;
12'h018:outb<=50'b00000000000000000000111111111111111111111111000000;
12'h019:outb<=50'b00000000000000000000000011111111111111000000000000;
12'h01a:outb<=50'b00000000000000000000000011111111111111000000000000;
12'h01b:outb<=50'b00000000000000000000000000000000000000000000000000;
12'h01c:outb<=50'b00000000000000000000000000000000000000000000000000;
12'h01d:outb<=50'b00000000000000000000000000000000000000000000000000;
12'h01e:outb<=50'b00000000000000000000000000000000000000000000000000;
12'h01f:outb<=50'b00000000000000000000000000000000000000000000000000;
12'h020:outb<=50'b00000000000000000000000000000000000000000000000000;
12'h021:outb<=50'b00000000000000000000000000000000000000000000000000;
12'h022:outb<=50'b00000000000000000000000000000000000000000000000000;
12'h023:outb<=50'b00000000000000000000000000000000000000000000000000;
12'h024:outb<=50'b00000000000000000000000000000000000000000000000000;
12'h025:outb<=50'b00000000000000000000000000000000000000000000000000;
12'h026:outb<=50'b00000000000000000000000000000000000000000000000000;

12'h100:outb<=50'b00000000000000000000000000000000000000000000000000;
12'h101:outb<=50'b00000000000000000000000000000000000000000000000000;
12'h102:outb<=50'b00000000000000000000000000000000000000000000000000;
12'h103:outb<=50'b00000000000000000000000000000000000000000000000000;
12'h104:outb<=50'b00000000000000000000000000000000000000000000000000;
12'h105:outb<=50'b00000000000000000000000000000000000000000000000000;
12'h106:outb<=50'b00000000000000000000000000000000000000000000000000;
12'h107:outb<=50'b00000000000000000000000000000000000000000000000000;
12'h108:outb<=50'b00000000000000000000000000000000000000000000000000;
12'h109:outb<=50'b00000000000000000000000000000000000000000000000000;
12'h10a:outb<=50'b00000000000000000000000000000000000000000000000000;
12'h10b:outb<=50'b00000000000011110000000000000000000000000000000000;
12'h10c:outb<=50'b00000000000011110000000000000000000000000000000000;
12'h10d:outb<=50'b00000000001111111100000000000000000000000000000000;
12'h10e:outb<=50'b00000000001111111100000000000000000000000000000000;
12'h10f:outb<=50'b00000000111111111111000000000000000000000000000000;
12'h100:outb<=50'b00000001111111111111000000000000000000000000000000;
12'h111:outb<=50'b00000011111111111111000000000000000000000000000000;
12'h112:outb<=50'b00000111111111111111000000000000000000000000000000;
12'h113:outb<=50'b00001111111111111111111111111111111111111111110000;
12'h114:outb<=50'b00001111111111111111111111111111111111111111110000;
12'h115:outb<=50'b00000000000000001111111111111111111111110000000000;
12'h116:outb<=50'b00000000000000001111111111111111111111110000000000;
12'h117:outb<=50'b00000000000000000000111111111111111111111111000000;
12'h118:outb<=50'b00000000000000000000111111111111111111111111000000;
12'h119:outb<=50'b00000000000000000000001111111111111100000000000000;
12'h11a:outb<=50'b00000000000000000000001111111111111100000000000000;
12'h11b:outb<=50'b00000000000000000000001111111111111000000000000000;
12'h11c:outb<=50'b00000000000000000000001111111111110000000000000000;
12'h11d:outb<=50'b00000000000000000000001111111111100000000000000000;
12'h11e:outb<=50'b00000000000000000000001111111111000000000000000000;
12'h11f:outb<=50'b00000000000000000000001111111110000000000000000000;
12'h120:outb<=50'b00000000000000000000001111111100000000000000000000;
12'h121:outb<=50'b00000000000000000000001111111000000000000000000000;
12'h122:outb<=50'b00000000000000000000001111110000000000000000000000;
12'h123:outb<=50'b00000000000000000000001111100000000000000000000000;
12'h124:outb<=50'b00000000000000000000001111000000000000000000000000;
12'h125:outb<=50'b00000000000000000000001110000000000000000000000000;
12'h126:outb<=50'b00000000000000000000001100000000000000000000000000;
endcase
end
endmodule

