module scorename_rom(vc,datas);
input [10:0] vc;
output reg [46:0] datas;
always@(vc)
        case((vc-7'd100))
4'd0:datas<=47'b00000000000000000000000000000000000000000000;
4'd1:datas<=47'b00000000000000000000000000000000000000000000;
4'd2:datas<=47'b11111110011111110000111000011111110011111110;
4'd3:datas<=47'b11111110011111110001101100011111110011111110;
4'd4:datas<=47'b11000000011000000011000110011000110011000000;
4'd5:datas<=47'b11000000011000000011000110011000110011000000;
4'd6:datas<=47'b11111110011000000011000110011111100011111110;
4'd7:datas<=47'b11111110011000000011000110011111100011111110;
4'd8:datas<=47'b00000110011000000011000110011000110011000000;
4'd9:datas<=47'b00000110011000000011000110011000110011000000;
4'd10:datas<=47'b11111110011111110001101100011000110011111110;
4'd11:datas<=47'b11111110011111110000111000011000110011111110;
4'd12:datas<=47'b00000000000000000000000000000000000000000000;
4'd13:datas<=47'b00000000000000000000000000000000000000000000;
4'd14:datas<=47'b00000000000000000000000000000000000000000000;
4'd15:datas<=47'b00000000000000000000000000000000000000000000;     
        endcase
endmodule