module gameover_rom(vc,outg);
input[10:0]vc;
output reg [249:0]outg;
always@(vc)
begin
case(vc-150)
7'd0:outg<=250'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000;
7'd1:outg<=250'b0000000000000000000000011111111111111100000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000011111111111111000000000000000000000000000000111111111111100000000000000000000000000000000000000011111111111111000000;
7'd2:outg<=250'b0000000000000000000111111111111111111111110011111100000000000000000000000000000000000111111111111100000000000000000000000000000000111111111111111111110000000000000000000000000011111111111111111000000111111111111111111111111111111111111111111111100000;
7'd3:outg<=250'b0000000000000000011111111111111111111111111111111110000000000000000000000000000000001111111111111110000000000000000000000000000001111111111111111111110000000000000000000000001111111111111111111100001111111111111111111111111111111111111111111111110000;
7'd4:outg<=250'b0000000000000001111111111111111111111111111111111111000000000000000000000000000000011111111111111111000000000000000000000000000011111111111111111111111000000000000000000000001111111111111111111110001111111111111111111111111111111111111111111111110000;
7'd5:outg<=250'b0000000000000111111111111111111111111111111111111111100000000000000000000000000000011111111111111111100000000000000000000000000011111111111111111111111000000000000000000000011111111111111111111110001111111111111111111111111111111111111111111111110000;
7'd6:outg<=250'b0000000000001111111111111111111111111111111111111111100000000000000000000000000000011111111111111111110000000000000000000000000011111111111111111111111100000000000000000000111111111111111111111110001111111111111111111111111111111111111111111111111000;
7'd7:outg<=250'b0000000000011111111111111111111111111111111111111111110000000000000000000000000000111111111111111111110000000000000000000000000011111111111111111111111100000000000000000000111111111111111111111110001111111111111111111111111111111111111111111111111000;
7'd8:outg<=250'b0000000001111111111111111111111111111111111111111111110000000000000000000000000000111111111111111111111000000000000000000000000001111111111111111111111110000000000000000000111111111111111111111100000001111111111111111111111111111111111111111111111000;
7'd9:outg<=250'b0000000011111111111111111111111111111111111111111111110000000000000000000000000000111111111111111111111100000000000000000000000000011111111111111111111111000000000000000001111111111111111111110000000000111111111111111111110000000000001111111111111000;
7'd10:outg<=250'b0000000011111111111111111111100000111111111111111111111000000000000000000000000000111111111111111111111100000000000000000000000000000111111111111111111111000000000000000001111111111111111111110000000000011111111111111111100000000000000001111111111000;
7'd11:outg<=250'b0000000111111111111111111100000000000111111111111111111000000000000000000000000000111111111111111111111110000000000000000000000000000111111111111111111111100000000000000011111111111111111111100000000000011111111111111111100000000000000000111111111000;
7'd12:outg<=250'b0000001111111111111111111000000000000011111111111111111000000000000000000000000000111111111111111111111110000000000000000000000000000011111111111111111111100000000000000111111111111111111111100000000000011111111111111111100000000000000000011111111000;
7'd13:outg<=250'b0000011111111111111111110000000000000000111111111111111000000000000000000000000000111111111111111111111111000000000000000000000000000011111111111111111111110000000000000111111111111111111111100000000000011111111111111111100000000000000000001111111000;
7'd14:outg<=250'b0000011111111111111111100000000000000000011111111111111000000000000000000000000000111111111111111111111111100000000000000000000000000011111111111111111111110000000000001111111111111111111111100000000000001111111111111111100000000000000000001111110000;
7'd15:outg<=250'b0000111111111111111111000000000000000000001111111111110000000000000000000000000000111111111111111111111111100000000000000000000000000011111111111111111111111000000000001111111111111111111111000000000000001111111111111111100000000011110000000111100000;
7'd16:outg<=250'b0000111111111111111111000000000000000000001111111111110000000000000000000000000001111111111111111111111111110000000000000000000000000011111111111111111111111000000000011111111111111111111111000000000000001111111111111111100000000111111000000000000000;
7'd17:outg<=250'b0001111111111111111110000000000000000000000111111111110000000000000000000000000001111111111111111111111111110000000000000000000000000011111111111111111111111100000000011111111111111111111111000000000000001111111111111111100000000111111000000000000000;
7'd18:outg<=250'b0001111111111111111110000000000000000000000011111111100000000000000000000000000001111111111111111111111111111000000000000000000000000011111111111111111111111100000000111111111111111111111111000000000000001111111111111111000000000111111100000000000000;
7'd19:outg<=250'b0011111111111111111110000000000000000000000000111110000000000000000000000000000011111111111111111111111111111000000000000000000000000011111111111111111111111110000000111111111111111111111111000000000000001111111111111111000000000111111100000000000000;
7'd20:outg<=250'b0011111111111111111110000000000000000000000000000000000000000000000000000000000011111111111111111111111111111100000000000000000000000011111111111111111111111111000001111111111111111111111111000000000000001111111111111111100000000111111100000000000000;
7'd21:outg<=250'b0011111111111111111110000000000000000000000000000000000000000000000000000000000111111111101111111111111111111100000000000000000000000011111111111111111111111111000001111111111111111111111111000000000000001111111111111111100000001111111100000000000000;
7'd22:outg<=250'b0011111111111111111100000000000000000000000000000000000000000000000000000000000111111111000111111111111111111110000000000000000000000011111111111111111111111111100011111111111111111111111111000000000000001111111111111111100000001111111100000000000000;
7'd23:outg<=250'b0111111111111111111100000000000000000000000000000000000000000000000000000000001111111110000011111111111111111110000000000000000000000011111111111111111111111111110111111111111111111111111111000000000000001111111111111111111111111111111110000000000000;
7'd24:outg<=250'b0111111111111111111110000000000000000000000000000000000000000000000000000000001111111110000001111111111111111111000000000000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111110000000000000;
7'd25:outg<=250'b0111111111111111111110000000000000000000000000000000000000000000000000000000011111111100000001111111111111111111000000000000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111110000000000000;
7'd26:outg<=250'b0111111111111111111110000000000000000000011111111110000000000000000000000000011111111100000000111111111111111111100000000000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111110000000000000;
7'd27:outg<=250'b0111111111111111111110000000000000001111111111111111111110000000000000000000011111111100000000111111111111111111100000000000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111110000000000000;
7'd28:outg<=250'b0111111111111111111110000000000001111111111111111111111111100000000000000000111111111000000000011111111111111111110000000000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111110000000000000;
7'd29:outg<=250'b0111111111111111111110000000000011111111111111111111111111110000000000000000111111111000000000011111111111111111110000000000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111110000000000000;
7'd30:outg<=250'b0111111111111111111110000000000111111111111111111111111111111000000000000001111111110000000000001111111111111111110000000000000000000011111111110011111111111111111111111111111111111111111111000000000000001111111111111111111001111111111100000000000000;
7'd31:outg<=250'b0111111111111111111111000000000111111111111111111111111111111000000000000001111111110000000000001111111111111111111000000000000000000011111111110001111111111111111111111100011111111111111111000000000000001111111111111111110000001111111100000000000000;
7'd32:outg<=250'b0011111111111111111111000000000111111111111111111111111111111000000000000011111111111000000000011111111111111111111000000000000000000011111111110001111111111111111111111000011111111111111111000000000000001111111111111111100000001111111100000000000000;
7'd33:outg<=250'b0011111111111111111111000000000111111111111111111111111111111000000000000011111111111111111111111111111111111111111100000000000000000011111111100000111111111111111111111000011111111111111111000000000000001111111111111111100000000111111100000000000000;
7'd34:outg<=250'b0011111111111111111111100000000011111111111111111111111111110000000000000111111111111111111111111111111111111111111100000000000000000011111111100000111111111111111111110000011111111111111111000000000000001111111111111111100000000111111000000000000000;
7'd35:outg<=250'b0011111111111111111111100000000000111111111111111111111111000000000000000111111111111111111111111111111111111111111110000000000000000011111111100000011111111111111111110000011111111111111111000000000000001111111111111111100000000111111000000000000000;
7'd36:outg<=250'b0001111111111111111111110000000000000011111111111111111100000000000000001111111111111111111111111111111111111111111110000000000000000011111111100000011111111111111111100000011111111111111111000000000000001111111111111111100000000111111000000000111110;
7'd37:outg<=250'b0001111111111111111111111000000000000001111111111111111000000000000000001111111111111111111111111111111111111111111111000000000000000011111111100000001111111111111111100000011111111111111111000000000000001111111111111111100000000011110000000000111111;
7'd38:outg<=250'b0000111111111111111111111000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111000000000000000111111111100000001111111111111111000000011111111111111111000000000000001111111111111111100000000000000000000001111111;
7'd39:outg<=250'b0000111111111111111111111100000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111100000000000000111111111100000001111111111111111000000011111111111111111000000000000001111111111111111100000000000000000000001111111;
7'd40:outg<=250'b0000011111111111111111111110000000000001111111111111110000000000000000111111111111111111111111111111111111111111111111100000000000000111111111100000000111111111111110000000011111111111111111000000000000001111111111111111100000000000000000000011111111;
7'd41:outg<=250'b0000011111111111111111111111000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111110000000000000111111111100000000111111111111110000000011111111111111111100000000000001111111111111111100000000000000000000111111111;
7'd42:outg<=250'b0000001111111111111111111111110000000111111111111111100000000000000001111111111110000000000000000011111111111111111111110000000000000111111111100000000011111111111100000000011111111111111111100000000000011111111111111111100000000000000000000111111111;
7'd43:outg<=250'b0000000111111111111111111111111111111111111111111111100000000000000001111111111100000000000000000000111111111111111111111000000000000111111111100000000011111111111100000000011111111111111111100000000000011111111111111111110000000000000000001111111111;
7'd44:outg<=250'b0000000111111111111111111111111111111111111111111111000000000000000011111111111100000000000000000000111111111111111111111000000000000111111111110000000001111111111100000000111111111111111111100000000000011111111111111111110000000000000000011111111111;
7'd45:outg<=250'b0000000011111111111111111111111111111111111111111110000000000000000111111111111100000000000000000000111111111111111111111100000000000111111111110000000001111111111000000000111111111111111111110000000000011111111111111111111000000000000001111111111110;
7'd46:outg<=250'b0000000001111111111111111111111111111111111111111110000000000000001111111111111111000000000000000001111111111111111111111111100000001111111111110000000000111111111000000001111111111111111111111000000000111111111111111111111111111111111111111111111110;
7'd47:outg<=250'b0000000000111111111111111111111111111111111111111100000000000001111111111111111111110000000000001111111111111111111111111111110000011111111111111100000000111111110000000011111111111111111111111100000001111111111111111111111111111111111111111111111110;
7'd48:outg<=250'b0000000000001111111111111111111111111111111111111000000000000011111111111111111111110000000000001111111111111111111111111111111001111111111111111110000000011111110000000111111111111111111111111110000111111111111111111111111111111111111111111111111100;
7'd49:outg<=250'b0000000000000111111111111111111111111111111111100000000000000011111111111111111111110000000000011111111111111111111111111111111011111111111111111111000000011111100000000111111111111111111111111110001111111111111111111111111111111111111111111111111100;
7'd50:outg<=250'b0000000000000001111111111111111111111111111111000000000000000011111111111111111111110000000000011111111111111111111111111111111011111111111111111111000000001111100000001111111111111111111111111110001111111111111111111111111111111111111111111111111000;
7'd51:outg<=250'b0000000000000000011111111111111111111111111100000000000000000011111111111111111111110000000000001111111111111111111111111111110011111111111111111111000000001111000000000111111111111111111111111110001111111111111111111111111111111111111111111111111000;
7'd52:outg<=250'b0000000000000000000111111111111111111111110000000000000000000011111111111111111111100000000000001111111111111111111111111111100011111111111111111110000000000110000000000111111111111111111111111100001111111111111111111111111111111111111111111111110000;
7'd53:outg<=250'b0000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000011111111111111111111111110000000111111111111111100000000000000000000000001111111111111111111110000000011111111111111111111111111111111111111111111100000;
7'd54:outg<=250'b0000000000000000000000000001111111000000000000000000000000000000000001111111100000000000000000000000000001111111111111000000000000000011111110000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000011000000;
7'd55:outg<=250'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd56:outg<=250'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd57:outg<=250'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd58:outg<=250'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd60:outg<=250'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd61:outg<=250'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd62:outg<=250'b0000000000000000000000001111111111110000000000000000000000000000000001111111111111111000000000000000000000011111111111111000000000000000000000000000000000000000001111111111000000000000001111100000000000001111111111111100000000000000000000000000000000;
7'd63:outg<=250'b0000000000000000000011111111111111111111000000000000000000000000011111111111111111111111100000000000000011111111111111111110000111111111111111111111111111111111111111111111000000000011111111111111111111111111111111111111100000000000000000000000000000;
7'd64:outg<=250'b0000000000000000011111111111111111111111110000000000000000000001111111111111111111111111111000000000001111111111111111111111001111111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111000000000000000000000000000;
7'd65:outg<=250'b0000000000000001111111111111111111111111111100000000000000000011111111111111111111111111111000000000011111111111111111111111011111111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111110000000000000000000000000;
7'd66:outg<=250'b0000000000000011111111111111111111111111111111000000000000000111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111000000000000000000000000;
7'd67:outg<=250'b0000000000001111111111111111111111111111111111110000000000000111111111111111111111111111111100000000011111111111111111111111011111111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111110000000000000000000000;
7'd68:outg<=250'b0000000000011111111111111111111111111111111111111000000000000111111111111111111111111111111000000000001111111111111111111111001111111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111110000000000000000000000;
7'd69:outg<=250'b0000000001111111111111111111111111111111111111111100000000000111111111111111111111111111110000000000000111111111111111111110000111111111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111000000000000000000000;
7'd70:outg<=250'b0000000001111111111111111111111111111111111111111110000000000011111111111111111111111111100000000000000011111111111111000000000001111111111111111111111000000000111111111111111000000001111111111111111111111111111111111111111111111100000000000000000000;
7'd71:outg<=250'b0000000011111111111111111111111111111111111111111111000000000000111111111111111111111111000000000000000001111111111110000000000000111111111111111111100000000000000011111111111000000000111111111111111111110000011111111111111111111100000000000000000000;
7'd72:outg<=250'b0000000111111111111111111111111111111111111111111111100000000000001111111111111111111111000000000000000001111111111110000000000000011111111111111111000000000000000001111111111000000000011111111111111111100000001111111111111111111100000000000000000000;
7'd73:outg<=250'b0000001111111111111111111000111111111111111111111111100000000000000111111111111111111111000000000000000001111111111100000000000000011111111111111111000000000000000000111111111000000000011111111111111111100000000111111111111111111100000000000000000000;
7'd74:outg<=250'b0000011111111111111111100000001111111111111111111111110000000000000111111111111111111111100000000000000011111111111100000000000000011111111111111111000000000000000000011111111000000000011111111111111111100000000111111111111111111110000000000000000000;
7'd75:outg<=250'b0000011111111111111111000000000011111111111111111111111000000000000011111111111111111111100000000000000011111111111000000000000000011111111111111111000000000000000000001111110000000000011111111111111111100000000111111111111111111110000000000000000000;
7'd76:outg<=250'b0000111111111111111110000000000001111111111111111111111000000000000011111111111111111111110000000000000111111111111000000000000000011111111111111111000000000001100000001111100000000000011111111111111111100000000111111111111111111110000000000000000000;
7'd77:outg<=250'b0000111111111111111110000000000000111111111111111111111100000000000001111111111111111111110000000000000111111111110000000000000000011111111111111111000000000111110000000011000000000000011111111111111111100000000111111111111111111110000000000000000000;
7'd78:outg<=250'b0001111111111111111100000000000000111111111111111111111100000000000001111111111111111111111000000000001111111111110000000000000000001111111111111111000000000111111000000000000000000000011111111111111111100000000111111111111111111100000000000000000000;
7'd79:outg<=250'b0001111111111111111100000000000000011111111111111111111110000000000000111111111111111111111000000000001111111111100000000000000000001111111111111111000000001111111000000000000000000000011111111111111111100000000111111111111111111100000000000000000000;
7'd80:outg<=250'b0011111111111111111100000000000000011111111111111111111110000000000000111111111111111111111100000000011111111111100000000000000000001111111111111111000000001111111000000000000000000000011111111111111111100000000111111111111111111100000000000000000000;
7'd81:outg<=250'b0011111111111111111100000000000000001111111111111111111110000000000000011111111111111111111100000000011111111111000000000000000000001111111111111111000000001111111100000000000000000000011111111111111111100000000111111111111111111000000000000000000000;
7'd82:outg<=250'b0011111111111111111100000000000000001111111111111111111111000000000000011111111111111111111100000000111111111111000000000000000000001111111111111111000000001111111100000000000000000000011111111111111111100000001111111111111111111000000000000000000000;
7'd83:outg<=250'b0011111111111111111100000000000000000111111111111111111111000000000000001111111111111111111110000000111111111110000000000000000000001111111111111111100000001111111100000000000000000000011111111111111111100000011111111111111111110000000000000000000000;
7'd84:outg<=250'b0111111111111111111100000000000000000111111111111111111111000000000000001111111111111111111110000001111111111110000000000000000000001111111111111111111111111111111100000000000000000000011111111111111111111111111111111111111111100000000000000000000000;
7'd85:outg<=250'b0111111111111111111100000000000000000111111111111111111111100000000000000111111111111111111111000001111111111100000000000000000000001111111111111111111111111111111100000000000000000000011111111111111111111111111111111111111111000000000000000000000000;
7'd86:outg<=250'b0111111111111111111110000000000000000011111111111111111111100000000000000111111111111111111111000011111111111100000000000000000000001111111111111111111111111111111100000000000000000000011111111111111111111111111111111111111110000000000000000000000000;
7'd87:outg<=250'b0111111111111111111110000000000000000011111111111111111111100000000000000111111111111111111111110111111111111000000000000000000000001111111111111111111111111111111100000000000000000000011111111111111111111111111111111111111000000000000000000000000000;
7'd88:outg<=250'b0111111111111111111110000000000000000011111111111111111111100000000000000011111111111111111111111111111111111000000000000000000000001111111111111111111111111111111100000000000000000000011111111111111111111111111111111111111000000000000000000000000000;
7'd89:outg<=250'b0111111111111111111110000000000000000001111111111111111111100000000000000011111111111111111111111111111111110000000000000000000000001111111111111111111111111111111100000000000000000000011111111111111111111111111111111111111100000000000000000000000000;
7'd90:outg<=250'b0111111111111111111111000000000000000001111111111111111111100000000000000001111111111111111111111111111111110000000000000000000000001111111111111111111111111111111100000000000000000000011111111111111111111111111111111111111111000000000000000000000000;
7'd91:outg<=250'b0111111111111111111111000000000000000001111111111111111111100000000000000001111111111111111111111111111111100000000000000000000000001111111111111111111111111111111100000000000000000000011111111111111111111111111111111111111111110000000000000000000000;
7'd92:outg<=250'b0111111111111111111111000000000000000001111111111111111111100000000000000000111111111111111111111111111111100000000000000000000000001111111111111111110000111111111100000000000000000000011111111111111111111111111111111111111111111000000000000000000000;
7'd93:outg<=250'b0111111111111111111111100000000000000001111111111111111111100000000000000000111111111111111111111111111111000000000000000000000000001111111111111111100000001111111100000000000000000000011111111111111111110001111111111111111111111100000000000000000000;
7'd94:outg<=250'b0011111111111111111111100000000000000001111111111111111111000000000000000000011111111111111111111111111111000000000000000000000000001111111111111111100000001111111100000000000000000000011111111111111111100000011111111111111111111110000000000000000000;
7'd95:outg<=250'b0011111111111111111111110000000000000001111111111111111111000000000000000000011111111111111111111111111110000000000000000000000000001111111111111111100000000111111000000000000000000000011111111111111111100000001111111111111111111110000000000000000000;
7'd96:outg<=250'b0011111111111111111111110000000000000001111111111111111111000000000000000000001111111111111111111111111100000000000000000000000000001111111111111111100000000111111000000000000000000000011111111111111111100000001111111111111111111111000000000000000000;
7'd97:outg<=250'b0011111111111111111111111000000000000001111111111111111111000000000000000000001111111111111111111111111100000000000000000000000000001111111111111111100000000111110000000000011100000000011111111111111111100000000111111111111111111111000000000000000000;
7'd98:outg<=250'b0001111111111111111111111000000000000001111111111111111110000000000000000000000111111111111111111111111100000000000000000000000000001111111111111111100000000111110000000001111110000000011111111111111111100000000111111111111111111111100000000000000000;
7'd99:outg<=250'b0001111111111111111111111100000000000001111111111111111110000000000000000000000111111111111111111111111000000000000000000000000000001111111111111111100000000011000000000001111111000000011111111111111111100000000111111111111111111111100000000000000000;
7'd100:outg<=250'b0000111111111111111111111100000000000001111111111111111100000000000000000000000111111111111111111111111000000000000000000000000000011111111111111111100000000000000000000011111111000000011111111111111111100000000011111111111111111111100000000000000000;
7'd101:outg<=250'b0000111111111111111111111110000000000011111111111111111100000000000000000000000011111111111111111111110000000000000000000000000000011111111111111111100000000000000000000011111111000000011111111111111111100000000011111111111111111111100000000000000000;
7'd102:outg<=250'b0000011111111111111111111111000000000011111111111111111000000000000000000000000011111111111111111111100000000000000000000000000000011111111111111111100000000000000000000111111111000000011111111111111111100000000011111111111111111111100000000000000000;
7'd103:outg<=250'b0000011111111111111111111111100000000111111111111111111000000000000000000000000001111111111111111111100000000000000000000000000000011111111111111111100000000000000000000111111111000000011111111111111111100000000011111111111111111111110000000000000000;
7'd104:outg<=250'b0000001111111111111111111111111000011111111111111111110000000000000000000000000001111111111111111111000000000000000000000000000000011111111111111111100000000000000000001111111111000000011111111111111111100000000001111111111111111111110000000000000000;
7'd105:outg<=250'b0000000111111111111111111111111111111111111111111111100000000000000000000000000000111111111111111111000000000000000000000000000000011111111111111111100000000000000000011111111110000000111111111111111111110000000001111111111111111111110000000000000000;
7'd106:outg<=250'b0000000111111111111111111111111111111111111111111111000000000000000000000000000000111111111111111111000000000000000000000000000000111111111111111111110000000000000001111111111110000001111111111111111111110000000001111111111111111111110000000000000000;
7'd107:outg<=250'b0000000011111111111111111111111111111111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000111111111111111111111100000000011111111111111110000011111111111111111111111000000000111111111111111111111100000000000000;
7'd108:outg<=250'b0000000001111111111111111111111111111111111111111100000000000000000000000000000000011111111111111100000000000000000000000000000001111111111111111111111111111111111111111111111110000111111111111111111111111100000000111111111111111111111111000000000000;
7'd109:outg<=250'b0000000000011111111111111111111111111111111111111000000000000000000000000000000000001111111111111100000000000000000000000000000111111111111111111111111111111111111111111111111100001111111111111111111111111110000000111111111111111111111111100000000000;
7'd110:outg<=250'b0000000000001111111111111111111111111111111111110000000000000000000000000000000000001111111111111000000000000000000000000000001111111111111111111111111111111111111111111111111100001111111111111111111111111111000000011111111111111111111111100000000000;
7'd111:outg<=250'b0000000000000111111111111111111111111111111111000000000000000000000000000000000000000111111111111000000000000000000000000000001111111111111111111111111111111111111111111111111000001111111111111111111111111111000000011111111111111111111111100000000000;
7'd112:outg<=250'b0000000000000001111111111111111111111111111100000000000000000000000000000000000000000111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111000001111111111111111111111111111000000001111111111111111111111100000000000;
7'd113:outg<=250'b0000000000000000011111111111111111111111110000000000000000000000000000000000000000000011111111110000000000000000000000000000001111111111111111111111111111111111111111111111110000000111111111111111111111111110000000000111111111111111111111000000000000;
7'd114:outg<=250'b0000000000000000000011111111111111111110000000000000000000000000000000000000000000000011111111100000000000000000000000000000000111111111111111111111111111111111111111111111100000000001111111111111111111111100000000000011111111111111111110000000000000;
7'd115:outg<=250'b0000000000000000000000001111111111100000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000001111111111111111100000000000000000111111111111111100000000000000;
7'd116:outg<=250'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000;
endcase
end
endmodule