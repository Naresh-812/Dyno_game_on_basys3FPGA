module cloud_rom(vc,c,outc);
input[10:0]vc;
input[10:0]c;
output reg [69:0]outc;
always@(vc)
begin
case(vc-c)

7'd0:outc<=70'b0000000000000000000000000000000000000000000000000000000000000000000000;
7'd1:outc<=70'b0000000000000000000000000001111100000000000000000000000000000000000000;
7'd2:outc<=70'b0000000000000000000000011111111111110000000000000000000000000000000000;
7'd3:outc<=70'b0000000000000000000001111111111111111100000000000000000000000000000000;
7'd4:outc<=70'b0000000000000000000011111111101111111110000000000000000000000000000000;
7'd5:outc<=70'b0000000000000000001111110000000000111111100000000000000000000000000000;
7'd6:outc<=70'b0000000000000000011111000000000000000111110000000000000000000000000000;
7'd7:outc<=70'b0000000000000000011110000000000000000011110000000000000000000000000000;
7'd8:outc<=70'b0000000000000000111100000000000000000001111000000000000000000000000000;
7'd9:outc<=70'b0000000000000001111000000000000000000000111100000000000000000000000000;
7'd10:outc<=70'b0000000000000001110000000000000000000000011100000000000000000000000000;
7'd11:outc<=70'b0000000000000011110000000000000000000000011110000000000000000000000000;
7'd12:outc<=70'b0000000000000011100000000000000000000000001111111111100000000000000000;
7'd13:outc<=70'b0000000000000111100000000000000000000000001111111111111000000000000000;
7'd14:outc<=70'b0000000001111111100000000000000000000000001111111111111110000000000000;
7'd15:outc<=70'b0000000111111111000000000000000000000000000111000000111111000000000000;
7'd16:outc<=70'b0000011111111111000000000000000000000000000100000000001111100000000000;
7'd17:outc<=70'b0000111111000000000000000000000000000000000000000000000011110000000000;
7'd18:outc<=70'b0001111100000000000000000000000000000000000000000000000001111000000000;
7'd19:outc<=70'b0001111000000000000000000000000000000000000000000000000001111000000000;
7'd20:outc<=70'b0011110000000000000000000000000000000000000000000000000000111100000000;
7'd21:outc<=70'b0011100000000000000000000000000000000000000000000000000000111100000000;
7'd22:outc<=70'b0111100000000000000000000000000000000000000000000000000000011110000000;
7'd23:outc<=70'b0111000000000000000000000000000000000000000000000000000000011111100000;
7'd24:outc<=70'b0111000000000000000000000000000000000000000000000000000000011111111000;
7'd25:outc<=70'b0111000000000000000000000000000000000000000000000000000000000011111100;
7'd26:outc<=70'b0111000000000000000000000000000000000000000000000000000000000000111100;
7'd27:outc<=70'b0111000000000000000000000000000000000000000000000000000000000000011110;
7'd28:outc<=70'b0111000000000000000000000000000000000000000000000000000000000000001110;
7'd29:outc<=70'b0111100000000000000000000000000000000000000000000000000000000000001110;
7'd30:outc<=70'b0011100000000000000000000000000000000000000000000000000000000000001110;
7'd31:outc<=70'b0011110000000000000000000000000000000000000000000000000000000000001110;
7'd32:outc<=70'b0001111000000000000000000000000000000000000000000000000000000000011110;
7'd33:outc<=70'b0000111100000000000000000000000000000000000000000000000000000000011100;
7'd34:outc<=70'b0000111111100000000000000000000000000000000000000000000000000001111100;
7'd35:outc<=70'b0000001111111111111111111111111111111111111111111111111111111111111000;
7'd36:outc<=70'b0000000111111111111111111111111111111111111111111111111111111111110000;
7'd37:outc<=70'b0000000001111111111111111111111111111111111111111111111111111111000000;
7'd38:outc<=70'b0000000000000000000000000000000000000000000000000000000000000000000000;

endcase
end
endmodule
