module catcus_rom( 
	input wire [11:0] addr,
	output reg [39:0] outtr
	);
	
always@(addr)
case((addr))

/////////////////////////////////////////////////catcus 1/////////////////////////////////////////////////////////////////
12'h100 : outtr <= 40'b000111000000000000000000000000000000000;
12'h101 : outtr <= 40'b001111100000000000000000000000000000000;
12'h102 : outtr <= 40'b011111110000000000000000000000000000000;
12'h103 : outtr <= 40'b011111110000000000000000000000000000000;
12'h104 : outtr <= 40'b011111110000000000000000000000000000000;
12'h105 : outtr <= 40'b011111111000000000000000000000000000000;
12'h106 : outtr <= 40'b111111111000000000000000000000000000000;
12'h107 : outtr <= 40'b111111111000000000000000000000000000000;
12'h108 : outtr <= 40'b011111111000000000000000000000000000000;
12'h109 : outtr <= 40'b011111111000000011111100000000000000000;
12'h10a : outtr <= 40'b001111110000000111111100000000000000000;
12'h10b : outtr <= 40'b001111110010000111111110000000000000000;
12'h10c : outtr <= 40'b000111110111100111111000000110000000000;
12'h10d : outtr <= 40'b000001111111111011111101111100000000000;
12'h10e : outtr <= 40'b000000011111111111100011111111000000000;
12'h10f : outtr <= 40'b000000111111111110000111111111100000000;
12'h110 : outtr <= 40'b000000011111111100001111111111100000000;
12'h111 : outtr <= 40'b000000011111111100001111111111100000000;
12'h112 : outtr <= 40'b000000001111111100001111111111100000000;
12'h113 : outtr <= 40'b000000001111111000001111111111100000000;
12'h114 : outtr <= 40'b000000000111111000001111111111100000000;
12'h115 : outtr <= 40'b000111111111110000010111111111000000000;
12'h116 : outtr <= 40'b000111111111100000000111111111000000000;
12'h117 : outtr <= 40'b001111111111100000000111111110000000000;
12'h118 : outtr <= 40'b010111111111100000000011111110000000000;
12'h119 : outtr <= 40'b000111111111000000000011111100000000000;
12'h11a : outtr <= 40'b000011111111001111111011111000000000000;
12'h11b : outtr <= 40'b000001111110111111111111100000000000000;
12'h11c : outtr <= 40'b000000111110111111111110000000000000000;
12'h11d : outtr <= 40'b000000001111111111111110000000000000000;
12'h11e : outtr <= 40'b000000000011111111111110000000000000000;
12'h11f : outtr <= 40'b000000000011111111111110000000000000000;
12'h120 : outtr <= 40'b000000000001111111111110000000000000000;
12'h121 : outtr <= 40'b000000000001111111111110000000000000000;
12'h122 : outtr <= 40'b000000000001111111111100000000000000000;
12'h123 : outtr <= 40'b000000000110111111111000000000000000000;
12'h124 : outtr <= 40'b000000000000111111111000000000000000000;
12'h125 : outtr <= 40'b000000000000011111111000000000000000000;
12'h126 : outtr <= 40'b000000000000011111110000000000000000000;
12'h127 : outtr <= 40'b000000000000001111110000000000000000000;
12'h128 : outtr <= 40'b000000000111111111111110000000000000000;
12'h129 : outtr <= 40'b111111111111111111111110000011100000000;
12'h12a : outtr <= 40'b000000000111100001110000000000000000000;

/////////////////////////////////////////////////catcus 2/////////////////////////////////////////////////////////////////

12'h200:outtr<=40'b0000000000000000000000000000000000000000;
12'h201:outtr<=40'b0000001000000000000000000000000000000000;
12'h202:outtr<=40'b0000011100000000000000000000000000000000;
12'h203:outtr<=40'b0000011100000000000000000000000000000000;
12'h204:outtr<=40'b0000011100000000000000000000000000000000;
12'h205:outtr<=40'b0000011100000000000000000000000000000000;
12'h206:outtr<=40'b0100011100000000000000000000000000000000;
12'h207:outtr<=40'b0110011100000000000000000000000000000000;
12'h208:outtr<=40'b0110011100000000000000000000000000000000;
12'h209:outtr<=40'b0110011100000000000000000000000000000000;
12'h20a:outtr<=40'b0110011100000000000000000000000000000000;
12'h20b:outtr<=40'b0110011100100000000000000000000000000000;
12'h20c:outtr<=40'b0110011100110000000000000000000000000000;
12'h20d:outtr<=40'b0110011100110000000000000000000000000000;
12'h20e:outtr<=40'b0110011100110000000000000000000000000000;
12'h20f:outtr<=40'b0110011100110000000000000000000000000000;
12'h210:outtr<=40'b0110011100110000000000000000000000000000;
12'h211:outtr<=40'b0110011100110000000000000000000000000000;
12'h212:outtr<=40'b0110011100110000000000000000000000000000;
12'h213:outtr<=40'b0110011100110000000000000000000000000000;
12'h214:outtr<=40'b0110011100110000000000000000000000000000;
12'h215:outtr<=40'b0111111100110000000000000000000000000000;
12'h216:outtr<=40'b0111111100110000000000000000000000000000;
12'h217:outtr<=40'b0011111100110000000000000000000000000000;
12'h218:outtr<=40'b0011111100110000000000000000000000000000;
12'h219:outtr<=40'b0001111100110000000000000000000000000000;
12'h21a:outtr<=40'b0000011100110000000000000000000000000000;
12'h21b:outtr<=40'b0000011111100000000000000000000000000000;
12'h21c:outtr<=40'b0000011111100000000000000000000000000000;
12'h21d:outtr<=40'b0000011111000000000000000000000000000000;
12'h22e:outtr<=40'b0000011111000000000000000000000000000000;
12'h22f:outtr<=40'b0000011100000000000000000000000000000000;
12'h220:outtr<=40'b0000011100000000000000000000000000000000;
12'h221:outtr<=40'b0000011100000000000000000000000000000000;
12'h222:outtr<=40'b0000011100000000000000000000000000000000;
12'h223:outtr<=40'b0000011100000000000000000000000000000000;
12'h224:outtr<=40'b0000011100000000000000000000000000000000;
12'h225:outtr<=40'b0000011100000000000000000000000000000000;
12'h226:outtr<=40'b0000011100000000000000000000000000000000;
12'h227:outtr<=40'b0000011100000000000000000000000000000000;
12'h228:outtr<=40'b0000011100000000000000000000000000000000;
12'h229:outtr<=40'b0000011100000000000000000000000000000000;
12'h22a:outtr<=40'b0000011100000000000000000000000000000000;

/////////////////////////////////////////////////catcus 3/////////////////////////////////////////////////////////////////

12'h300:outtr<=40'b0000000000000000001100000000000000000000;
12'h301:outtr<=40'b0000000000000000001110000000000000000000;
12'h302:outtr<=40'b0000100000000000001110000000000000000000;
12'h303:outtr<=40'b0000110000000000001110000000000000000000;
12'h304:outtr<=40'b0000110000000000001110000000000000000000;
12'h305:outtr<=40'b0000110000000000001110000000000000000000;
12'h306:outtr<=40'b0000110000000010001110000000000000000000;
12'h307:outtr<=40'b0000110000000011001110000000000000000000;
12'h308:outtr<=40'b0000110010000011001110000000000000000000;
12'h309:outtr<=40'b0000110010000011001110000000000000000000;
12'h30a:outtr<=40'b0000110010000011001110000000000000000000;
12'h30b:outtr<=40'b0000110010000011001110010000000000000000;
12'h30c:outtr<=40'b0000110010000011001110011000000000000000;
12'h30d:outtr<=40'b0000110010000011001110011000000000000000;
12'h30e:outtr<=40'b0000110010000011001110011000000000000000;
12'h30f:outtr<=40'b0000110010000011001110011000000000000000;
12'h310:outtr<=40'b0100110010000011001110011000000000000000;
12'h311:outtr<=40'b0100111110000011001110011000000000000000;
12'h312:outtr<=40'b0100111100000011001110011000000000000000;
12'h313:outtr<=40'b0100111100000011001110011000000000000000;
12'h314:outtr<=40'b0100110000100011111110011000000000000000;
12'h315:outtr<=40'b0100110000100011111110011000000000000000;
12'h316:outtr<=40'b0100110000100011111110011000000000000000;
12'h317:outtr<=40'b0100110000100001111110011000000000000000;
12'h318:outtr<=40'b0100110000100001111110011000000000000000;
12'h319:outtr<=40'b0100110010100100001110011000000000000000;
12'h31a:outtr<=40'b0100110010100100001110010000000000000000;
12'h31b:outtr<=40'b0100110010100100001111110000000000000000;
12'h31c:outtr<=40'b0100110010100100001111100000000000000000;
12'h31d:outtr<=40'b0111110010100100001111100000000000000000;
12'h31e:outtr<=40'b0111110010100100001110000000000000000000;
12'h31f:outtr<=40'b0011110010100100001110000000000000000000;
12'h320:outtr<=40'b0011110010100100001110000000000000000000;
12'h321:outtr<=40'b0000110010100100001110000000000000000000;
12'h322:outtr<=40'b0000110011111000001110000000000000000000;
12'h323:outtr<=40'b0000110001111000001110000000000000000000;
12'h324:outtr<=40'b0000110001100000001110000000000000000000;
12'h325:outtr<=40'b0000110000100000001110000000000000000000;
12'h326:outtr<=40'b0000110000100000001110000000000000000000;
12'h327:outtr<=40'b0000110000100000001110000000000000000000;
12'h328:outtr<=40'b0000110000100000001110000000000000000000;
12'h329:outtr<=40'b0000110000100000001110000000000000000000;
12'h32a:outtr<=40'b0000110000100000001110000000000000000000;


/////////////////////////////////////////////////catcus 4/////////////////////////////////////////////////////////////////

12'h400 : outtr <= 40'b000000000011111100000000000000000000000;
12'h401 : outtr <= 40'b000000000111111110000000000000000000000;
12'h402 : outtr <= 40'b000000000111111100000000000000000000000;
12'h403 : outtr <= 40'b000000000111111110000000000000000000000;
12'h404 : outtr <= 40'b000000000111111110000000000000000000000;
12'h405 : outtr <= 40'b000000000111111100000000000000000000000;
12'h406 : outtr <= 40'b000000000011111100000000000000000000000;
12'h407 : outtr <= 40'b000000000111111110000000000000000000000;
12'h408 : outtr <= 40'b000000000111111100000000000000000000000;
12'h409 : outtr <= 40'b000000001111111100000000000000000000000;
12'h40a : outtr <= 40'b000000000111111100011110000000000000000;
12'h40b : outtr <= 40'b000000001111111100111110000000000000000;
12'h40c : outtr <= 40'b000000000111111100111110000000000000000;
12'h40d : outtr <= 40'b000000000111111110011110000000000000000;
12'h40e : outtr <= 40'b000000000111111100111111000000000000000;
12'h40f : outtr <= 40'b011100000111111100011110000000000000000;
12'h410 : outtr <= 40'b111111000111111100111110000000000000000;
12'h411 : outtr <= 40'b111111000111111100111111000001111000000;
12'h412 : outtr <= 40'b111111001111111100111111000001111000000;
12'h413 : outtr <= 40'b111111100111111110111110000001111001110;
12'h414 : outtr <= 40'b111111000111111110111110000001111101110;
12'h415 : outtr <= 40'b111111000111111101111110000001111001100;
12'h416 : outtr <= 40'b111111000111111110111100000001111101100;
12'h417 : outtr <= 40'b111111000111111100111100110001111001100;
12'h418 : outtr <= 40'b111111000111111111111000111001111111100;
12'h419 : outtr <= 40'b111111001111111101110000111001111111000;
12'h41a : outtr <= 40'b111111000111111111100000111111111110011;
12'h41b : outtr <= 40'b111111100111111110000000111101111100111;
12'h41c : outtr <= 40'b111111000111111110000000011111111000111;
12'h41d : outtr <= 40'b011111101111111100000000001111111101111;
12'h41e : outtr <= 40'b011111100111111110000000001111111001110;
12'h41f : outtr <= 40'b001111110111111100000000000001111111110;
12'h420 : outtr <= 40'b000111111111111100000000000001111111100;
12'h421 : outtr <= 40'b000111111111111100000000000001111111000;
12'h422 : outtr <= 40'b000000111111111100000000000001111100000;
12'h423 : outtr <= 40'b000000000111111100000000000001111000000;
12'h424 : outtr <= 40'b000000000111111100000000000001111000000;
12'h425 : outtr <= 40'b000000000111111111000000000001111000000;
12'h426 : outtr <= 40'b000000000111111100000000000001111100000;
12'h427 : outtr <= 40'b000000000111111100000000000001111100000;
12'h428 : outtr <= 40'b000000000111111100000000000001111100000;
12'h429 : outtr <= 40'b000000000111111100000000000001111100000;
12'h42a : outtr <= 40'b000000000111111100000000000001111100000;

/////////////////////////////////////////////////catcus 5/////////////////////////////////////////////////////////////////
12'h500 : outtr <= 40'b000111000000000000000000000000000000000;
12'h501 : outtr <= 40'b001111100000000000000000000000000000000;
12'h502 : outtr <= 40'b011111110000000000000000000000000000000;
12'h503 : outtr <= 40'b011111110000000000000000000000000000000;
12'h504 : outtr <= 40'b011111110000000000000000000000000000000;
12'h505 : outtr <= 40'b011111111000000000000000000000000000000;
12'h506 : outtr <= 40'b111111111000000000000000000000000000000;
12'h507 : outtr <= 40'b111111111000000000000000000000000000000;
12'h508 : outtr <= 40'b011111111000000000000000000000000000000;
12'h509 : outtr <= 40'b011111111000000011111100000000000000000;
12'h50a : outtr <= 40'b001111110000000111111100000000000000000;
12'h50b : outtr <= 40'b001111110010000111111110000000000000000;
12'h50c : outtr <= 40'b000111110111100111111000000110000000000;
12'h50d : outtr <= 40'b000001111111111011111101111100000000000;
12'h50e : outtr <= 40'b000000011111111111100011111111000000000;
12'h50f : outtr <= 40'b000000111111111110000111111111100000000;
12'h510 : outtr <= 40'b000000011111111100001111111111100000000;
12'h511 : outtr <= 40'b000000011111111100001111111111100000000;
12'h512 : outtr <= 40'b000000001111111100001111111111100000000;
12'h513 : outtr <= 40'b000000001111111000001111111111100000000;
12'h514 : outtr <= 40'b000000000111111000001111111111100000000;
12'h515 : outtr <= 40'b000111111111110000010111111111000000000;
12'h516 : outtr <= 40'b000111111111100000000111111111000000000;
12'h517 : outtr <= 40'b001111111111100000000111111110000000000;
12'h518 : outtr <= 40'b010111111111100000000011111110000000000;
12'h519 : outtr <= 40'b000111111111000000000011111100000000000;
12'h51a : outtr <= 40'b000011111111001111111011111000000000000;
12'h51b : outtr <= 40'b000001111110111111111111100000000000000;
12'h51c : outtr <= 40'b000000111110111111111110000000000000000;
12'h51d : outtr <= 40'b000000001111111111111110000000000000000;
12'h51e : outtr <= 40'b000000000011111111111110000000000000000;
12'h51f : outtr <= 40'b000000000011111111111110000000000000000;
12'h520 : outtr <= 40'b000000000001111111111110000000000000000;
12'h521 : outtr <= 40'b000000000001111111111110000000000000000;
12'h522 : outtr <= 40'b000000000001111111111100000000000000000;
12'h523 : outtr <= 40'b000000000110111111111000000000000000000;
12'h524 : outtr <= 40'b000000000000111111111000000000000000000;
12'h525 : outtr <= 40'b000000000000011111111000000000000000000;
12'h526 : outtr <= 40'b000000000000011111110000000000000000000;
12'h527 : outtr <= 40'b000000000000001111110000000000000000000;
12'h528 : outtr <= 40'b000000000111111111111110000000000000000;
12'h529 : outtr <= 40'b111111111111111111111110000011100000000;
12'h52a : outtr <= 40'b000000000111100001110000000000000000000;
default: outtr <= 40'b0;

endcase
endmodule
