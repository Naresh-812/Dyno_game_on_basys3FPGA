module dinodown_rom(vc,outdd);
input [10:0]vc;
output reg [49:0]outdd;
always@(vc)
begin
case(vc-11'd374)
5'd0:outdd<=50'b00000000000000000000000000000000000000000000000000;
5'd1:outdd<=50'b00000000000000000000000000000000000000000000000000;
5'd2:outdd<=50'b00000000000000000000000000000000000000000000000000;
5'd3:outdd<=50'b00000000000000000000000000000000000000000000000000;
5'd4:outdd<=50'b00000000000000000000000000000000000000000000000000;
5'd5:outdd<=50'b00000000000000000000000000000000000000000000000000;
5'd6:outdd<=50'b00000000000000000000000000000000000000000000000000;
5'd7:outdd<=50'b00010000000000000000000000000000000000000000000000;
5'd8:outdd<=50'b00011000000000000000000000000000011111111111110000;
5'd9:outdd<=50'b00011111000000111111111111110001111111111111111000;
5'd10:outdd<=50'b00011111111111111111111111111111110011111111111000;
5'd11:outdd<=50'b00001111111111111111111111111111110011111111111000;
5'd12:outdd<=50'b00000111111111111111111111111111111111111111111000;
5'd13:outdd<=50'b00000011111111111111111111111111111111111111111000;
5'd14:outdd<=50'b00000011111111111111111111111111111111111111111000;
5'd15:outdd<=50'b00000000111111111111111111111111111111111111111000;
5'd16:outdd<=50'b00000000011111111111111111111111111111100000000000;
5'd17:outdd<=50'b00000000011111111111111111111111111111100000000000;
5'd18:outdd<=50'b00000000000111111111111111111000011111111111000000;
5'd19:outdd<=50'b00000000000011111111111111111000000000000000000000;
5'd20:outdd<=50'b00000000000001111111110000110000000000000000000000;
5'd21:outdd<=50'b00000000000011110000111100110000000000000000000000;
5'd22:outdd<=50'b00000000000011100000000000111000000000000000000000;
5'd23:outdd<=50'b00000000000011100000000000000000000000000000000000;
5'd24:outdd<=50'b00000000000010000000000000000000000000000000000000;
5'd25:outdd<=50'b00000000000010000000000000000000000000000000000000;
5'd26:outdd<=50'b00000000000011100000000000000000000000000000000000;
5'd27:outdd<=50'b00000000000000000000000000000000000000000000000000;
5'd28:outdd<=50'b00000000000000000000000000000000000000000000000000;
endcase
end
endmodule